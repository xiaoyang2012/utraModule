// megafunction wizard: %ALTOCT%VBB%
// GENERATION: STANDARD
// VERSION: WM1.0
// MODULE: ALT_OCT_POWER 

// ============================================================
// File Name: DDR3_OCT.v
// Megafunction Name(s):
// 			ALT_OCT_POWER
//
// Simulation Library Files(s):
// 			altera_mf
// ============================================================
// ************************************************************
// THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
//
// 12.1 Build 177 11/07/2012 SJ Full Version
// ************************************************************

//Copyright (C) 1991-2012 Altera Corporation
//Your use of Altera Corporation's design tools, logic functions 
//and other software and tools, and its AMPP partner logic 
//functions, and any output files from any of the foregoing 
//(including device programming or simulation files), and any 
//associated documentation or information are expressly subject 
//to the terms and conditions of the Altera Program License 
//Subscription Agreement, Altera MegaCore Function License 
//Agreement, or other applicable license agreement, including, 
//without limitation, that your use is for the sole purpose of 
//programming logic devices manufactured by Altera and sold by 
//Altera or its authorized distributors.  Please refer to the 
//applicable agreement for further details.

module DDR3_OCT (
	rzqin,
	parallelterminationcontrol,
	seriesterminationcontrol)/* synthesis synthesis_clearbox = 1 */;

	input	[0:0]  rzqin;
	output	[15:0]  parallelterminationcontrol;
	output	[15:0]  seriesterminationcontrol;

endmodule

// ============================================================
// CNX file retrieval info
// ============================================================
// Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Cyclone V"
// Retrieval info: PRIVATE: SYNTH_WRAPPER_GEN_POSTFIX STRING "0"
// Retrieval info: CONSTANT: INTENDED_DEVICE_FAMILY STRING "Cyclone V"
// Retrieval info: CONSTANT: LPM_TYPE STRING "ALT_OCT_POWER"
// Retrieval info: CONSTANT: width_ptc NUMERIC "16"
// Retrieval info: CONSTANT: width_stc NUMERIC "16"
// Retrieval info: USED_PORT: parallelterminationcontrol 0 0 16 0 OUTPUT NODEFVAL "parallelterminationcontrol[15..0]"
// Retrieval info: USED_PORT: rzqin 0 0 1 0 INPUT NODEFVAL "rzqin[0..0]"
// Retrieval info: USED_PORT: seriesterminationcontrol 0 0 16 0 OUTPUT NODEFVAL "seriesterminationcontrol[15..0]"
// Retrieval info: CONNECT: @rzqin 0 0 1 0 rzqin 0 0 1 0
// Retrieval info: CONNECT: parallelterminationcontrol 0 0 16 0 @parallelterminationcontrol 0 0 16 0
// Retrieval info: CONNECT: seriesterminationcontrol 0 0 16 0 @seriesterminationcontrol 0 0 16 0
// Retrieval info: GEN_FILE: TYPE_NORMAL DDR3_OCT.v TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL DDR3_OCT.inc FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL DDR3_OCT.cmp FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL DDR3_OCT.bsf FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL DDR3_OCT_inst.v FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL DDR3_OCT_bb.v TRUE
// Retrieval info: LIB_FILE: altera_mf
